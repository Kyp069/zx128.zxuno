//-------------------------------------------------------------------------------------------------
module audio
//-------------------------------------------------------------------------------------------------
(
	input  wire      clock,
	input  wire      reset,
	input  wire[7:0] specdrum,
	input  wire      speaker,
	input  wire      mic,
	input  wire      ear,
	input  wire[7:0] a1,
	input  wire[7:0] b1,
	input  wire[7:0] c1,
	input  wire[7:0] a2,
	input  wire[7:0] b2,
	input  wire[7:0] c2,
	output wire[1:0] audio
);
//-------------------------------------------------------------------------------------------------

wire[2:0] sem = { speaker, ear, mic };

wire[7:0] ula
	= sem == 3'b000 ? 8'h00
	: sem == 3'b001 ? 8'h24
	: sem == 3'b010 ? 8'h40
	: sem == 3'b011 ? 8'h64
	: sem == 3'b100 ? 8'hB8
	: sem == 3'b101 ? 8'hC0
	: sem == 3'b110 ? 8'hF8
	:     /* 3'b111 */8'hFF;

//-------------------------------------------------------------------------------------------------

reg[3:0] cc;
always @(posedge clock) if(cc == 8) cc <= 1'd0; else cc <= cc+1'd1;

wire[7:0] l;
wire[7:0] r;

assign { l, r }
	= cc == 0 ? { 2{ula} }
	: cc == 1 ? { a1, c1 }
	: cc == 2 ? { a1, c1 }
	: cc == 3 ? { 2{b1} }
	: cc == 4 ? { a2, c2 }
	: cc == 5 ? { a2, c2 }
	: cc == 6 ? { 2{b2} }
	: cc == 7 ? { 2{specdrum} }
	: /* == 8 */{ 2{specdrum} };

//-------------------------------------------------------------------------------------------------

dac #(.MSBI(7)) L
(
	.clock  (clock  ),
	.reset  (reset  ),
	.d      (l      ),
	.q      (audio[0])
);

dac #(.MSBI(7)) R
(
	.clock  (clock  ),
	.reset  (reset  ),
	.d      (r      ),
	.q      (audio[1])
);

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
