//-------------------------------------------------------------------------------------------------
module dpr
//-------------------------------------------------------------------------------------------------
#
(
	parameter AW = 14
)
(
	input  wire         clock,
	input  wire         ce1,
	input  wire         we1,
	input  wire[   7:0] d1,
	input  wire[AW-1:0] a1,
	input  wire         ce2,
	output reg [   7:0] q2,
	input  wire[AW-1:0] a2
);
//-------------------------------------------------------------------------------------------------

reg[7:0] ram[(2**AW)-1:0];

always @(posedge clock) if(ce1) if(!we1) ram[a1] <= d1;
always @(posedge clock) if(ce2) q2 <= ram[a2];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
